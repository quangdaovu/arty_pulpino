
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [10:0]  A,
    output logic [31:0] Q
  );

  const logic [0:1099] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hEF410113,
    32'h00001D17,
    32'hF5CD0D13,
    32'h00001D97,
    32'hF58D8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h688000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h46811101,
    32'h45A14601,
    32'hCE064515,
    32'h7C0000EF,
    32'h02000513,
    32'h015000EF,
    32'h45014581,
    32'h045000EF,
    32'h02000593,
    32'h00EF0028,
    32'h00EF0FF0,
    32'h55330670,
    32'h3CE31005,
    32'h4681FE15,
    32'h45A14601,
    32'h07000513,
    32'h78C000EF,
    32'h02000513,
    32'h7E0000EF,
    32'h45014581,
    32'h011000EF,
    32'h02000593,
    32'h00EF0068,
    32'h00EF0CB0,
    32'h55330330,
    32'h3CE31005,
    32'h2703FE15,
    32'h37B300C1,
    32'hE789F077,
    32'h00814503,
    32'h00A03533,
    32'h01C12083,
    32'h80826105,
    32'h45A11101,
    32'h46014681,
    32'hCE064519,
    32'hCA26CC22,
    32'hC64EC84A,
    32'h734000EF,
    32'h00EF4501,
    32'h458178A0,
    32'h00EF4505,
    32'h00EF7BA0,
    32'h54337E60,
    32'h3CE31005,
    32'h46A1FE14,
    32'h061385B6,
    32'h051305F0,
    32'h00EF0610,
    32'h450170A0,
    32'h760000EF,
    32'h85224581,
    32'h790000EF,
    32'h7BC000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h00009537,
    32'h051345D5,
    32'h00EFC7C5,
    32'h00EF10F0,
    32'h45811B30,
    32'h00EF4521,
    32'h043771A0,
    32'h09B700FF,
    32'h6905FF01,
    32'h00FF84B7,
    32'h00841613,
    32'h02000693,
    32'h051345A1,
    32'h00EF0EB0,
    32'h65216B60,
    32'h70C000EF,
    32'h45094581,
    32'h73C000EF,
    32'h01340533,
    32'h944A65A1,
    32'h7F4000EF,
    32'hFC941AE3,
    32'h758000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h00009537,
    32'h051345B5,
    32'h00EFC945,
    32'h00EF0AB0,
    32'h458114F0,
    32'h00EF4521,
    32'h89B76B60,
    32'h6905FF10,
    32'h010004B7,
    32'h00841613,
    32'h02000693,
    32'h051345A1,
    32'h00EF0EB0,
    32'h65216560,
    32'h6AC000EF,
    32'h45094581,
    32'h6DC000EF,
    32'h01340533,
    32'h944A65A1,
    32'h794000EF,
    32'hFC941AE3,
    32'h00009537,
    32'h02200593,
    32'hCA450513,
    32'h055000EF,
    32'h0F9000EF,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000313,
    32'h208367A5,
    32'h240301C1,
    32'h24830181,
    32'h29030141,
    32'h29830101,
    32'hA82300C1,
    32'h61050667,
    32'h71398302,
    32'hD452DC22,
    32'h4A376461,
    32'hDA26000F,
    32'hD05AD256,
    32'hCC62CE5E,
    32'hD84ADE06,
    32'hCA66D64E,
    32'hC66EC86A,
    32'h00009C37,
    32'h00009BB7,
    32'h00009B37,
    32'h00009AB7,
    32'h240A0A13,
    32'h000094B7,
    32'h6A040413,
    32'h468145A1,
    32'h05134601,
    32'h00EF0660,
    32'h45015AE0,
    32'h604000EF,
    32'h45054581,
    32'h634000EF,
    32'h660000EF,
    32'h10055933,
    32'hFE193CE3,
    32'h468145A1,
    32'h05134601,
    32'h00EF0990,
    32'h45015860,
    32'h5DC000EF,
    32'h854A4581,
    32'h60C000EF,
    32'h638000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h468145A1,
    32'h05134601,
    32'h00EF0660,
    32'h450155E0,
    32'h5B4000EF,
    32'h450D4581,
    32'h5E4000EF,
    32'h610000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h468145A1,
    32'h05134601,
    32'h00EF0990,
    32'h45015360,
    32'h58C000EF,
    32'h450D4581,
    32'h5BC000EF,
    32'h5E8000EF,
    32'h10055933,
    32'hFE193CE3,
    32'h000097B7,
    32'hCC878513,
    32'h00EF45B5,
    32'h45A173A0,
    32'h46014681,
    32'h00EF4519,
    32'h45015020,
    32'h558000EF,
    32'h854A4581,
    32'h588000EF,
    32'h5B4000EF,
    32'h10055933,
    32'hFE193CE3,
    32'h46E145A1,
    32'hFF000637,
    32'h0D800513,
    32'h4D8000EF,
    32'h00EF4501,
    32'h458152E0,
    32'h00EF854A,
    32'h00EF55E0,
    32'h553358A0,
    32'h3CE31005,
    32'hF0EFFE15,
    32'hC519CEFF,
    32'h00EF8552,
    32'hF0EF79E0,
    32'hF97DCE3F,
    32'h000097B7,
    32'hCA078513,
    32'h00EF4585,
    32'h97B76CA0,
    32'h05930000,
    32'h851302E0,
    32'h00EFCD87,
    32'h09376BA0,
    32'h00EF00FF,
    32'h0DB775A0,
    32'h4D37FF01,
    32'h45A100FF,
    32'h46014681,
    32'h00EF4519,
    32'h45014720,
    32'h4C8000EF,
    32'h45054581,
    32'h01B909B3,
    32'h4F4000EF,
    32'h520000EF,
    32'h10055CB3,
    32'hFE1CBCE3,
    32'h161346E1,
    32'h45A10089,
    32'h00EF4509,
    32'h05134460,
    32'h00EF4000,
    32'h458149A0,
    32'h00EF8566,
    32'h05934CA0,
    32'h854E4000,
    32'h50C000EF,
    32'h4EC000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h08090913,
    32'h8513A811,
    32'h00EFD084,
    32'h00EF63E0,
    32'h85226E20,
    32'h6F4000EF,
    32'hC39FF0EF,
    32'hF5654585,
    32'hF9A911E3,
    32'h000097B7,
    32'hD0C78513,
    32'h00EF4589,
    32'h97B761A0,
    32'h05930000,
    32'h85130290,
    32'h00EFD107,
    32'h893760A0,
    32'h00EF00FF,
    32'h8DB76AA0,
    32'hCD37FF10,
    32'h45A100FF,
    32'h46014681,
    32'h00EF4519,
    32'h45013C20,
    32'h418000EF,
    32'h45054581,
    32'h01B909B3,
    32'h444000EF,
    32'h470000EF,
    32'h10055CB3,
    32'hFE1CBCE3,
    32'h161346E1,
    32'h45A10089,
    32'h00EF4509,
    32'h05133960,
    32'h00EF4000,
    32'h45813EA0,
    32'h00EF8566,
    32'h059341A0,
    32'h854E4000,
    32'h45C000EF,
    32'h43C000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h08090913,
    32'h8513A811,
    32'h00EFD084,
    32'h00EF58E0,
    32'h85226320,
    32'h644000EF,
    32'hB89FF0EF,
    32'hF5654585,
    32'hF9A911E3,
    32'h000097B7,
    32'h85134599,
    32'h00EFD387,
    32'h099356A0,
    32'h00EF0310,
    32'h091360A0,
    32'h0D130320,
    32'hA0290330,
    32'h09250D63,
    32'hD7A506E3,
    32'h03D00593,
    32'hD40C0513,
    32'h544000EF,
    32'h5E8000EF,
    32'h02800593,
    32'hD80B8513,
    32'h534000EF,
    32'h5D8000EF,
    32'h02700593,
    32'hDACB0513,
    32'h524000EF,
    32'h5C8000EF,
    32'h02C00593,
    32'hDD4A8513,
    32'h514000EF,
    32'h5B8000EF,
    32'h558000EF,
    32'hFB351AE3,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000313,
    32'h208367A5,
    32'h240303C1,
    32'h24830381,
    32'h29030341,
    32'h29830301,
    32'h2A0302C1,
    32'h2A830281,
    32'h2B030241,
    32'h2B830201,
    32'h2C0301C1,
    32'h2C830181,
    32'h2D030141,
    32'h2D830101,
    32'hA82300C1,
    32'h61210667,
    32'h20838302,
    32'h240303C1,
    32'h24830381,
    32'h29030341,
    32'h29830301,
    32'h2A0302C1,
    32'h2A830281,
    32'h2B030241,
    32'h2B830201,
    32'h2C0301C1,
    32'h2C830181,
    32'h2D030141,
    32'h2D830101,
    32'h612100C1,
    32'hB11FF06F,
    32'hCC221101,
    32'hC84ACA26,
    32'hC452C64E,
    32'hC05AC256,
    32'h9A37CE06,
    32'h99B70000,
    32'h99370000,
    32'h94B70000,
    32'h04130000,
    32'h0A930310,
    32'h0B130320,
    32'hA0290330,
    32'h09550263,
    32'h0B650263,
    32'h03D00593,
    32'hD40A0513,
    32'h440000EF,
    32'h4E4000EF,
    32'h02800593,
    32'hD8098513,
    32'h430000EF,
    32'h4D4000EF,
    32'h02700593,
    32'hDAC90513,
    32'h420000EF,
    32'h4C4000EF,
    32'h02C00593,
    32'hDD448513,
    32'h410000EF,
    32'h4B4000EF,
    32'h454000EF,
    32'hFA851AE3,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000313,
    32'h4B0267A5,
    32'h01C12083,
    32'h01812403,
    32'h01412483,
    32'h01012903,
    32'h00C12983,
    32'h00812A03,
    32'h00412A83,
    32'h0667A823,
    32'h83026105,
    32'h20834B02,
    32'h240301C1,
    32'h24830181,
    32'h29030141,
    32'h29830101,
    32'h2A0300C1,
    32'h2A830081,
    32'h61050041,
    32'hA39FF06F,
    32'h20834B02,
    32'h240301C1,
    32'h24830181,
    32'h29030141,
    32'h29830101,
    32'h2A0300C1,
    32'h2A830081,
    32'h61050041,
    32'hB67FF06F,
    32'h45051101,
    32'hCC22CE06,
    32'hC84ACA26,
    32'hC452C64E,
    32'h00EFC256,
    32'h45E90AA0,
    32'h00EF4501,
    32'h94B730E0,
    32'h47110098,
    32'h1A1027B7,
    32'hC3D86925,
    32'h8493440D,
    32'h9AB76804,
    32'h99B70000,
    32'h09130000,
    32'h9A37E3C9,
    32'h85260000,
    32'h3B0000EF,
    32'h02B00593,
    32'h8513E531,
    32'hC839E049,
    32'h330000EF,
    32'h00890533,
    32'h00EF4585,
    32'h45A13260,
    32'hE30A0513,
    32'h31C000EF,
    32'h3C0000EF,
    32'h38E3147D,
    32'h2083FDF4,
    32'h450101C1,
    32'h01812403,
    32'h01412483,
    32'h01012903,
    32'h00C12983,
    32'h00812A03,
    32'h00412A83,
    32'h80826105,
    32'h85134585,
    32'h00EFCA0A,
    32'hF0EF2E60,
    32'hB7E9E63F,
    32'h00009537,
    32'h05134585,
    32'h00EFCA05,
    32'hF0EF2D20,
    32'hBF7595BF,
    32'hFF010113,
    32'h00812423,
    32'h00000593,
    32'h00050413,
    32'h00F00513,
    32'h00112623,
    32'h39C000EF,
    32'h00000593,
    32'h00E00513,
    32'h390000EF,
    32'h00000593,
    32'h00D00513,
    32'h384000EF,
    32'h00000593,
    32'h00C00513,
    32'h378000EF,
    32'h04805663,
    32'h00000593,
    32'h01000513,
    32'h368000EF,
    32'h02142E63,
    32'h00000593,
    32'h00B00513,
    32'h358000EF,
    32'h02242663,
    32'h00000593,
    32'h00000513,
    32'h348000EF,
    32'h00342E63,
    32'h00C12083,
    32'h00812403,
    32'h00000593,
    32'h00100513,
    32'h01010113,
    32'h32C0006F,
    32'h00C12083,
    32'h00812403,
    32'h01010113,
    32'h00008067,
    32'h00004837,
    32'hF0080813,
    32'h00869693,
    32'h02000713,
    32'h1A1027B7,
    32'h40B70733,
    32'h0106F6B3,
    32'hF265B5B3,
    32'h00E51533,
    32'h00878813,
    32'h00C78713,
    32'h00B6E5B3,
    32'h01078793,
    32'h00A82023,
    32'h00C72023,
    32'h00B7A023,
    32'h00008067,
    32'h01059593,
    32'h10055533,
    32'h00A5E5B3,
    32'h1A1027B7,
    32'h00B7AA23,
    32'h00008067,
    32'h1A102737,
    32'h01070713,
    32'h00072783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12783,
    32'h1007D7B3,
    32'h01051513,
    32'h00F56533,
    32'h00A12623,
    32'h00C12783,
    32'h00F72023,
    32'h01010113,
    32'h00008067,
    32'h00100793,
    32'h00858593,
    32'h00B795B3,
    32'h00A79533,
    32'h000017B7,
    32'hF0078793,
    32'h00F5F5B3,
    32'hEE853533,
    32'h00A5E533,
    32'h1A1027B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A1027B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'hD45597B3,
    32'hFF010113,
    32'hF455B5B3,
    32'h00F12423,
    32'h00058863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h00012623,
    32'h00C12603,
    32'h1A102737,
    32'h00812783,
    32'h00700693,
    32'h01870593,
    32'h02F65C63,
    32'h00072783,
    32'h0187D793,
    32'hFEF6ECE3,
    32'h00C12783,
    32'h00279793,
    32'h20F57783,
    32'h00F5A023,
    32'h00C12783,
    32'h00178793,
    32'h00F12623,
    32'h00C12603,
    32'h00812783,
    32'hFCF648E3,
    32'h01010113,
    32'h00008067,
    32'hD45597B3,
    32'hFF010113,
    32'hF455B5B3,
    32'h00F12423,
    32'h00058863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h00012623,
    32'h00C12683,
    32'h1A102737,
    32'h00812783,
    32'h02070813,
    32'h02F6DE63,
    32'h00072783,
    32'hCF0797B3,
    32'hFE078CE3,
    32'h00C12783,
    32'h00082583,
    32'h00C12683,
    32'h00168693,
    32'h00D12623,
    32'h01010613,
    32'h00279793,
    32'hFFC62603,
    32'h00812683,
    32'h00B567A3,
    32'hFCD646E3,
    32'h01010113,
    32'h00008067,
    32'h1A107737,
    32'h00470713,
    32'h00072603,
    32'h1A1007B7,
    32'hC0164633,
    32'h00C72023,
    32'h00478693,
    32'h00C78513,
    32'h0085D813,
    32'h08300713,
    32'h0FF5F593,
    32'h00E52023,
    32'h0106A023,
    32'h0A700713,
    32'h00B7A42B,
    32'h00E7A023,
    32'h00300793,
    32'h00F52023,
    32'h0006A783,
    32'h0F07F793,
    32'hC017C7B3,
    32'h00F6A023,
    32'h00008067,
    32'h04058263,
    32'h1A100637,
    32'h01460813,
    32'h00082783,
    32'h0207F793,
    32'hFE078CE3,
    32'h00150713,
    32'h0405468B,
    32'h1A1007B7,
    32'h00D7A023,
    32'hFFF58593,
    32'h03F450FB,
    32'h00058C63,
    32'h0017468B,
    32'hFFF58593,
    32'h00D62023,
    32'hFC0596E3,
    32'h00008067,
    32'h00008067,
    32'h1A100737,
    32'h01470713,
    32'h00072783,
    32'hFC17B7B3,
    32'hFE078CE3,
    32'h1A1007B7,
    32'h0007A503,
    32'h0FF57513,
    32'h00008067,
    32'h1A100737,
    32'h01472783,
    32'hFC17B7B3,
    32'h00078863,
    32'h00072503,
    32'h0FF57513,
    32'h00008067,
    32'hFF010113,
    32'h00112623,
    32'h02C000EF,
    32'h00C12083,
    32'h00000513,
    32'h01010113,
    32'h00008067,
    32'h1A100737,
    32'h01470713,
    32'h00072783,
    32'h0407F793,
    32'hFE078CE3,
    32'h00008067,
    32'hFF010113,
    32'h00A12623,
    32'h00C12783,
    32'h00F05C63,
    32'h00000793,
    32'h00000013,
    32'h00178793,
    32'h00C12703,
    32'hFEE7CAE3,
    32'h01010113,
    32'h00008067,
    32'h1A1076B7,
    32'h0006A783,
    32'hFF010113,
    32'h00F12623,
    32'h00100793,
    32'h00A797B3,
    32'h00C12703,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h00F12623,
    32'h00C12783,
    32'h00A595B3,
    32'h00F5E533,
    32'h00A12623,
    32'h00C12783,
    32'h00F6A023,
    32'h01010113,
    32'h00008067,
    32'h79706F43,
    32'h20676E69,
    32'h74736E49,
    32'h74637572,
    32'h736E6F69,
    32'h0000000A,
    32'h79706F43,
    32'h20676E69,
    32'h61746144,
    32'h0000000A,
    32'h656E6F44,
    32'h756A202C,
    32'h6E69706D,
    32'h6F742067,
    32'h736E4920,
    32'h63757274,
    32'h6E6F6974,
    32'h4D415220,
    32'h00000A2E,
    32'h61656C43,
    32'h656D2072,
    32'h79726F6D,
    32'h0000000A,
    32'h74697257,
    32'h6E492065,
    32'h75727473,
    32'h6F697463,
    32'h654D206E,
    32'h79726F6D,
    32'h6E6F6320,
    32'h746E6574,
    32'h206F7420,
    32'h20495053,
    32'h73616C66,
    32'h00000A68,
    32'h0000002E,
    32'h00000A0A,
    32'h74697257,
    32'h61442065,
    32'h4D206174,
    32'h726F6D65,
    32'h6F632079,
    32'h6E65746E,
    32'h6F742074,
    32'h49505320,
    32'h616C6620,
    32'h000A6873,
    32'h656E6F44,
    32'h00000A21,
    32'h65725020,
    32'h31207373,
    32'h206F7420,
    32'h72617473,
    32'h78652074,
    32'h74756365,
    32'h206E6F69,
    32'h6D6F7266,
    32'h61747320,
    32'h6F207472,
    32'h6E492066,
    32'h75727473,
    32'h6F697463,
    32'h656D206E,
    32'h79726F6D,
    32'h0000000A,
    32'h65725020,
    32'h32207373,
    32'h206F7420,
    32'h79706F63,
    32'h6F727020,
    32'h6D617267,
    32'h6F726620,
    32'h5053206D,
    32'h6C662049,
    32'h0A687361,
    32'h00000000,
    32'h65725020,
    32'h33207373,
    32'h206F7420,
    32'h74697277,
    32'h72702065,
    32'h6172676F,
    32'h6F74206D,
    32'h49505320,
    32'h616C6620,
    32'h000A6873,
    32'h20724F20,
    32'h73657270,
    32'h6E612073,
    32'h79656B79,
    32'h206F7420,
    32'h70736964,
    32'h2079616C,
    32'h73696874,
    32'h6E656D20,
    32'h67612075,
    32'h0A6E6961,
    32'h00000000,
    32'h7475410D,
    32'h6F62206F,
    32'h6620746F,
    32'h206D6F72,
    32'h20495053,
    32'h73616C46,
    32'h69772068,
    32'h73206C6C,
    32'h74726174,
    32'h74666120,
    32'h00207265,
    32'h63657320,
    32'h73646E6F,
    32'h00000000,
    32'h33323130,
    32'h37363534,
    32'h42413938,
    32'h46454443,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000014,
    32'h00000018,
    32'hFFFFF2E8,
    32'h00000084,
    32'h200E4200,
    32'h7F01114A,
    32'h00000020,
    32'h00000030,
    32'hFFFFF354,
    32'h00000152,
    32'h200E4200,
    32'h7F011152,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h0000003C,
    32'h00000054,
    32'hFFFFF482,
    32'h000003A2,
    32'h400E4200,
    32'h7E081144,
    32'h5C7A1411,
    32'h117D0911,
    32'h16117915,
    32'h77171178,
    32'h11761811,
    32'h12117F01,
    32'h7B13117C,
    32'h11751911,
    32'h1B11741A,
    32'h00000073,
    32'h0000002C,
    32'h00000094,
    32'hFFFFF7E4,
    32'h000000FC,
    32'h200E4200,
    32'h7E081150,
    32'h117D0911,
    32'h13117C12,
    32'h7A14117B,
    32'h11791511,
    32'h01117816,
    32'h0000007F,
    32'h00000028,
    32'h000000C4,
    32'hFFFFF8B0,
    32'h000000BC,
    32'h200E4200,
    32'h7F011150,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h00007915,
    32'h00000018,
    32'h000000F0,
    32'hFFFFF940,
    32'h0000009C,
    32'h100E4400,
    32'h7E081148,
    32'h7F01114C,
    32'h00000010,
    32'h0000010C,
    32'hFFFFF9C0,
    32'h00000044,
    32'h00000000,
    32'h00000010,
    32'h00000120,
    32'hFFFFF9F0,
    32'h00000018,
    32'h00000000,
    32'h00000010,
    32'h00000134,
    32'hFFFFF9F4,
    32'h00000038,
    32'h100E5000,
    32'h00000010,
    32'h00000148,
    32'hFFFFFA18,
    32'h00000030,
    32'h00000000,
    32'h00000010,
    32'h0000015C,
    32'hFFFFFA34,
    32'h0000001C,
    32'h100E4C00,
    32'h00000010,
    32'h00000170,
    32'hFFFFFA3C,
    32'h00000078,
    32'h100E4800,
    32'h00000010,
    32'h00000184,
    32'hFFFFFAA0,
    32'h00000078,
    32'h100E4800,
    32'h00000010,
    32'h00000198,
    32'hFFFFFB04,
    32'h0000005C,
    32'h00000000,
    32'h00000010,
    32'h000001AC,
    32'hFFFFFB4C,
    32'h0000004C,
    32'h00000000,
    32'h00000010,
    32'h000001C0,
    32'hFFFFFB84,
    32'h00000024,
    32'h00000000,
    32'h00000014,
    32'h000001D4,
    32'hFFFFFB94,
    32'h00000038,
    32'h100E6000,
    32'h7F011144,
    32'h00000010,
    32'h000001EC,
    32'hFFFFFBB4,
    32'h00000018,
    32'h00000000,
    32'h00000010,
    32'h00000200,
    32'hFFFFFBB8,
    32'h0000002C,
    32'h100E4400,
    32'h00000010,
    32'h00000214,
    32'hFFFFFBD0,
    32'h00000048,
    32'h100E4C00,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [10:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule